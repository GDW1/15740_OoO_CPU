module test ();

    initial begin
        $display("Test");
    end
endmodule
